-------------------------------------------------------------------------------
-- Title      : user_driver_pkg
-- Project    : DTP2
-------------------------------------------------------------------------------
-- File       : user_driver_pkg.vhd
-- Author     : Hans-Joachim Gelke
-- Company    : 
-- Created    : 2018-10-21
-- Last update: 2019-2-13
-- Platform   : 
-- Standard   : VHDL'08
-------------------------------------------------------------------------------
-- Description: For Students to add their own drivers
-------------------------------------------------------------------------------
-- Copyright (c) 2018 - 2019
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-02-13  1.0      Hans-Joachim    Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use work.simulation_pkg.all;

package user_driver_pkg is





end user_driver_pkg;

package body user_driver_pkg is



 

end user_driver_pkg;
