brudi@PAVEL-LAPTOP.13156:1620044363