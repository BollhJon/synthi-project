library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package reg_controller_pkg is    -- untested...

    type t_reg_array is array (0 to 5) of std_logic_vector(3 downto 0);

end package;
